--------------------------------------------------------------------------------
----                                                                        ----
---- Copyright (c) 2009, Sandro Amato                                       ----
---- All rights reserved.                                                   ----
----                                                                        ----
---- Redistribution  and  use in  source  and binary forms, with or without ----
---- modification,  are  permitted  provided that  the following conditions ----
---- are met:                                                               ----
----                                                                        ----
----     * Redistributions  of  source  code  must  retain the above        ----
----       copyright   notice,  this  list  of  conditions  and  the        ----
----       following disclaimer.                                            ----
----     * Redistributions  in  binary form must reproduce the above        ----
----       copyright   notice,  this  list  of  conditions  and  the        ----
----       following  disclaimer in  the documentation and/or  other        ----
----       materials provided with the distribution.                        ----
----     * Neither  the  name  of  SANDRO AMATO nor the names of its        ----
----       contributors may be used to  endorse or  promote products        ----
----       derived from this software without specific prior written        ----
----       permission.                                                      ----
----                                                                        ----
---- THIS SOFTWARE IS PROVIDED  BY THE COPYRIGHT  HOLDERS AND  CONTRIBUTORS ----
---- "AS IS"  AND  ANY EXPRESS OR  IMPLIED  WARRANTIES, INCLUDING,  BUT NOT ----
---- LIMITED  TO, THE  IMPLIED  WARRANTIES  OF MERCHANTABILITY  AND FITNESS ----
---- FOR  A PARTICULAR  PURPOSE  ARE  DISCLAIMED. IN  NO  EVENT  SHALL  THE ----
---- COPYRIGHT  OWNER  OR CONTRIBUTORS  BE LIABLE FOR ANY DIRECT, INDIRECT, ----
---- INCIDENTAL,  SPECIAL,  EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, ----
---- BUT  NOT LIMITED  TO,  PROCUREMENT OF  SUBSTITUTE  GOODS  OR SERVICES; ----
---- LOSS  OF  USE,  DATA,  OR PROFITS;  OR  BUSINESS INTERRUPTION) HOWEVER ----
---- CAUSED  AND  ON  ANY THEORY  OF LIABILITY, WHETHER IN CONTRACT, STRICT ----
---- LIABILITY,  OR  TORT  (INCLUDING  NEGLIGENCE  OR OTHERWISE) ARISING IN ----
---- ANY  WAY OUT  OF THE  USE  OF  THIS  SOFTWARE,  EVEN IF ADVISED OF THE ----
---- POSSIBILITY OF SUCH DAMAGE.                                            ----
--------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;


--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity charmaps_ROM is
  port (
    i_EN    : in  std_logic;            -- RAM Enable Input
    i_clock : in  std_logic;            -- Clock
    i_ADDR  : in  std_logic_vector (10 downto 0);  -- 11-bit Address Input
    o_DO    : out std_logic_vector(7 downto 0)  -- 8-bit Data Output
    );
end charmaps_ROM;

architecture Behavioral of charmaps_ROM is
  signal s_EN : std_logic;
  
  constant c_rom_size : natural := 2**11;

  type t_rom is array (c_rom_size-1 downto 0) of
    std_logic_vector (7 downto 0);

  constant c_rom : t_rom := (
    -- AUTOMATICALLY GENERATED... START

    0 => X"00", 1 => X"00", 2 => X"00", 3 => X"00", 
    4 => X"00", 5 => X"00", 6 => X"00", 7 => X"00", 
    8 => X"00", 9 => X"00", 10 => X"00", 11 => X"00", 
    12 => X"00", 13 => X"00", 14 => X"00", 15 => X"00", 
    16 => X"00", 17 => X"00", 18 => X"00", 19 => X"FF", 
    20 => X"00", 21 => X"00", 22 => X"FF", 23 => X"00", 
    24 => X"00", 25 => X"FF", 26 => X"00", 27 => X"00", 
    28 => X"FF", 29 => X"00", 30 => X"00", 31 => X"00", 
    32 => X"00", 33 => X"00", 34 => X"FF", 35 => X"00", 
    36 => X"00", 37 => X"FF", 38 => X"00", 39 => X"00", 
    40 => X"FF", 41 => X"00", 42 => X"00", 43 => X"FF", 
    44 => X"00", 45 => X"00", 46 => X"00", 47 => X"00", 
    48 => X"00", 49 => X"00", 50 => X"24", 51 => X"24", 
    52 => X"24", 53 => X"24", 54 => X"24", 55 => X"24", 
    56 => X"24", 57 => X"24", 58 => X"24", 59 => X"24", 
    60 => X"24", 61 => X"24", 62 => X"00", 63 => X"00", 
    64 => X"00", 65 => X"00", 66 => X"49", 67 => X"49", 
    68 => X"49", 69 => X"49", 70 => X"49", 71 => X"49", 
    72 => X"49", 73 => X"49", 74 => X"49", 75 => X"49", 
    76 => X"49", 77 => X"49", 78 => X"00", 79 => X"00", 
    80 => X"00", 81 => X"00", 82 => X"92", 83 => X"92", 
    84 => X"92", 85 => X"92", 86 => X"92", 87 => X"92", 
    88 => X"92", 89 => X"92", 90 => X"92", 91 => X"92", 
    92 => X"92", 93 => X"92", 94 => X"00", 95 => X"00", 
    96 => X"00", 97 => X"00", 98 => X"55", 99 => X"55", 
    100 => X"55", 101 => X"55", 102 => X"55", 103 => X"55", 
    104 => X"55", 105 => X"55", 106 => X"55", 107 => X"55", 
    108 => X"55", 109 => X"55", 110 => X"00", 111 => X"00", 
    112 => X"00", 113 => X"00", 114 => X"AA", 115 => X"AA", 
    116 => X"AA", 117 => X"AA", 118 => X"AA", 119 => X"AA", 
    120 => X"AA", 121 => X"AA", 122 => X"AA", 123 => X"AA", 
    124 => X"AA", 125 => X"AA", 126 => X"00", 127 => X"00", 
    128 => X"00", 129 => X"00", 130 => X"00", 131 => X"FF", 
    132 => X"00", 133 => X"FF", 134 => X"00", 135 => X"FF", 
    136 => X"00", 137 => X"FF", 138 => X"00", 139 => X"FF", 
    140 => X"00", 141 => X"FF", 142 => X"00", 143 => X"00", 
    144 => X"00", 145 => X"00", 146 => X"FC", 147 => X"F3", 
    148 => X"FC", 149 => X"F3", 150 => X"FC", 151 => X"F3", 
    152 => X"FC", 153 => X"F3", 154 => X"FC", 155 => X"F3", 
    156 => X"FC", 157 => X"F3", 158 => X"00", 159 => X"00", 
    160 => X"00", 161 => X"00", 162 => X"3F", 163 => X"CF", 
    164 => X"3F", 165 => X"CF", 166 => X"3F", 167 => X"CF", 
    168 => X"3F", 169 => X"CF", 170 => X"3F", 171 => X"CF", 
    172 => X"3F", 173 => X"CF", 174 => X"00", 175 => X"00", 
    176 => X"00", 177 => X"00", 178 => X"03", 179 => X"0C", 
    180 => X"03", 181 => X"0C", 182 => X"03", 183 => X"0C", 
    184 => X"03", 185 => X"0C", 186 => X"03", 187 => X"0C", 
    188 => X"03", 189 => X"0C", 190 => X"00", 191 => X"00", 
    192 => X"00", 193 => X"00", 194 => X"C0", 195 => X"30", 
    196 => X"C0", 197 => X"30", 198 => X"C0", 199 => X"30", 
    200 => X"C0", 201 => X"30", 202 => X"C0", 203 => X"30", 
    204 => X"C0", 205 => X"30", 206 => X"00", 207 => X"00", 
    208 => X"00", 209 => X"00", 210 => X"00", 211 => X"66", 
    212 => X"66", 213 => X"66", 214 => X"66", 215 => X"00", 
    216 => X"00", 217 => X"66", 218 => X"66", 219 => X"66", 
    220 => X"66", 221 => X"00", 222 => X"00", 223 => X"00", 
    224 => X"00", 225 => X"00", 226 => X"FF", 227 => X"99", 
    228 => X"99", 229 => X"99", 230 => X"99", 231 => X"FF", 
    232 => X"FF", 233 => X"99", 234 => X"99", 235 => X"99", 
    236 => X"99", 237 => X"FF", 238 => X"00", 239 => X"00", 
    240 => X"00", 241 => X"00", 242 => X"0F", 243 => X"0F", 
    244 => X"0F", 245 => X"0F", 246 => X"0F", 247 => X"0F", 
    248 => X"0F", 249 => X"0F", 250 => X"0F", 251 => X"0F", 
    252 => X"0F", 253 => X"0F", 254 => X"00", 255 => X"00", 
    256 => X"00", 257 => X"00", 258 => X"F0", 259 => X"F0", 
    260 => X"F0", 261 => X"F0", 262 => X"F0", 263 => X"F0", 
    264 => X"F0", 265 => X"F0", 266 => X"F0", 267 => X"F0", 
    268 => X"F0", 269 => X"F0", 270 => X"00", 271 => X"00", 
    272 => X"00", 273 => X"00", 274 => X"FF", 275 => X"FF", 
    276 => X"FF", 277 => X"FF", 278 => X"FF", 279 => X"FF", 
    280 => X"00", 281 => X"00", 282 => X"00", 283 => X"00", 
    284 => X"00", 285 => X"00", 286 => X"00", 287 => X"00", 
    288 => X"00", 289 => X"00", 290 => X"00", 291 => X"00", 
    292 => X"00", 293 => X"00", 294 => X"00", 295 => X"00", 
    296 => X"FF", 297 => X"FF", 298 => X"FF", 299 => X"FF", 
    300 => X"FF", 301 => X"FF", 302 => X"00", 303 => X"00", 
    304 => X"00", 305 => X"00", 306 => X"0F", 307 => X"0F", 
    308 => X"0F", 309 => X"0F", 310 => X"0F", 311 => X"0F", 
    312 => X"0F", 313 => X"0F", 314 => X"0F", 315 => X"0F", 
    316 => X"0F", 317 => X"0F", 318 => X"00", 319 => X"00", 
    320 => X"00", 321 => X"00", 322 => X"F0", 323 => X"F0", 
    324 => X"F0", 325 => X"F0", 326 => X"F0", 327 => X"F0", 
    328 => X"F0", 329 => X"F0", 330 => X"F0", 331 => X"F0", 
    332 => X"F0", 333 => X"F0", 334 => X"00", 335 => X"00", 
    336 => X"00", 337 => X"00", 338 => X"00", 339 => X"7E", 
    340 => X"42", 341 => X"42", 342 => X"42", 343 => X"42", 
    344 => X"42", 345 => X"42", 346 => X"42", 347 => X"42", 
    348 => X"7E", 349 => X"00", 350 => X"00", 351 => X"00", 
    352 => X"00", 353 => X"00", 354 => X"FF", 355 => X"81", 
    356 => X"81", 357 => X"81", 358 => X"81", 359 => X"81", 
    360 => X"81", 361 => X"81", 362 => X"81", 363 => X"81", 
    364 => X"81", 365 => X"FF", 366 => X"00", 367 => X"00", 
    368 => X"00", 369 => X"00", 370 => X"49", 371 => X"24", 
    372 => X"49", 373 => X"24", 374 => X"49", 375 => X"24", 
    376 => X"49", 377 => X"24", 378 => X"49", 379 => X"24", 
    380 => X"49", 381 => X"24", 382 => X"00", 383 => X"00", 
    384 => X"00", 385 => X"00", 386 => X"92", 387 => X"24", 
    388 => X"92", 389 => X"24", 390 => X"92", 391 => X"24", 
    392 => X"92", 393 => X"24", 394 => X"92", 395 => X"24", 
    396 => X"92", 397 => X"24", 398 => X"00", 399 => X"00", 
    400 => X"00", 401 => X"00", 402 => X"92", 403 => X"49", 
    404 => X"92", 405 => X"49", 406 => X"92", 407 => X"49", 
    408 => X"92", 409 => X"49", 410 => X"92", 411 => X"49", 
    412 => X"92", 413 => X"49", 414 => X"00", 415 => X"00", 
    416 => X"00", 417 => X"00", 418 => X"AA", 419 => X"55", 
    420 => X"AA", 421 => X"55", 422 => X"AA", 423 => X"55", 
    424 => X"AA", 425 => X"55", 426 => X"AA", 427 => X"55", 
    428 => X"AA", 429 => X"55", 430 => X"00", 431 => X"00", 
    432 => X"00", 433 => X"00", 434 => X"55", 435 => X"AA", 
    436 => X"55", 437 => X"AA", 438 => X"55", 439 => X"AA", 
    440 => X"55", 441 => X"AA", 442 => X"55", 443 => X"AA", 
    444 => X"55", 445 => X"AA", 446 => X"00", 447 => X"00", 
    448 => X"00", 449 => X"00", 450 => X"B6", 451 => X"DB", 
    452 => X"B6", 453 => X"DB", 454 => X"B6", 455 => X"DB", 
    456 => X"B6", 457 => X"DB", 458 => X"B6", 459 => X"DB", 
    460 => X"B6", 461 => X"DB", 462 => X"00", 463 => X"00", 
    464 => X"00", 465 => X"00", 466 => X"6D", 467 => X"DB", 
    468 => X"6D", 469 => X"DB", 470 => X"6D", 471 => X"DB", 
    472 => X"6D", 473 => X"DB", 474 => X"6D", 475 => X"DB", 
    476 => X"6D", 477 => X"DB", 478 => X"00", 479 => X"00", 
    480 => X"00", 481 => X"00", 482 => X"6D", 483 => X"B6", 
    484 => X"6D", 485 => X"B6", 486 => X"6D", 487 => X"B6", 
    488 => X"6D", 489 => X"B6", 490 => X"6D", 491 => X"B6", 
    492 => X"6D", 493 => X"B6", 494 => X"00", 495 => X"00", 
    496 => X"00", 497 => X"00", 498 => X"FF", 499 => X"FF", 
    500 => X"FF", 501 => X"FF", 502 => X"FF", 503 => X"FF", 
    504 => X"FF", 505 => X"FF", 506 => X"FF", 507 => X"FF", 
    508 => X"FF", 509 => X"FF", 510 => X"00", 511 => X"00", 
    512 => X"00", 513 => X"00", 514 => X"00", 515 => X"00", 
    516 => X"00", 517 => X"00", 518 => X"00", 519 => X"00", 
    520 => X"00", 521 => X"00", 522 => X"00", 523 => X"00", 
    524 => X"00", 525 => X"00", 526 => X"00", 527 => X"00", 
    528 => X"00", 529 => X"00", 530 => X"10", 531 => X"10", 
    532 => X"10", 533 => X"10", 534 => X"10", 535 => X"10", 
    536 => X"10", 537 => X"10", 538 => X"00", 539 => X"00", 
    540 => X"10", 541 => X"00", 542 => X"00", 543 => X"00", 
    544 => X"00", 545 => X"00", 546 => X"44", 547 => X"44", 
    548 => X"44", 549 => X"44", 550 => X"44", 551 => X"00", 
    552 => X"00", 553 => X"00", 554 => X"00", 555 => X"00", 
    556 => X"00", 557 => X"00", 558 => X"00", 559 => X"00", 
    560 => X"00", 561 => X"00", 562 => X"44", 563 => X"44", 
    564 => X"FE", 565 => X"44", 566 => X"44", 567 => X"44", 
    568 => X"44", 569 => X"44", 570 => X"FE", 571 => X"44", 
    572 => X"44", 573 => X"00", 574 => X"00", 575 => X"00", 
    576 => X"00", 577 => X"00", 578 => X"7C", 579 => X"92", 
    580 => X"90", 581 => X"90", 582 => X"90", 583 => X"7C", 
    584 => X"12", 585 => X"12", 586 => X"12", 587 => X"92", 
    588 => X"7C", 589 => X"00", 590 => X"00", 591 => X"00", 
    592 => X"00", 593 => X"00", 594 => X"60", 595 => X"90", 
    596 => X"92", 597 => X"64", 598 => X"08", 599 => X"10", 
    600 => X"20", 601 => X"4C", 602 => X"92", 603 => X"12", 
    604 => X"0C", 605 => X"00", 606 => X"00", 607 => X"00", 
    608 => X"00", 609 => X"00", 610 => X"30", 611 => X"48", 
    612 => X"88", 613 => X"88", 614 => X"90", 615 => X"70", 
    616 => X"50", 617 => X"8A", 618 => X"84", 619 => X"84", 
    620 => X"7A", 621 => X"00", 622 => X"00", 623 => X"00", 
    624 => X"00", 625 => X"00", 626 => X"10", 627 => X"10", 
    628 => X"10", 629 => X"10", 630 => X"10", 631 => X"00", 
    632 => X"00", 633 => X"00", 634 => X"00", 635 => X"00", 
    636 => X"00", 637 => X"00", 638 => X"00", 639 => X"00", 
    640 => X"00", 641 => X"00", 642 => X"10", 643 => X"20", 
    644 => X"20", 645 => X"40", 646 => X"40", 647 => X"40", 
    648 => X"40", 649 => X"40", 650 => X"20", 651 => X"20", 
    652 => X"10", 653 => X"00", 654 => X"00", 655 => X"00", 
    656 => X"00", 657 => X"00", 658 => X"10", 659 => X"08", 
    660 => X"08", 661 => X"04", 662 => X"04", 663 => X"04", 
    664 => X"04", 665 => X"04", 666 => X"08", 667 => X"08", 
    668 => X"10", 669 => X"00", 670 => X"00", 671 => X"00", 
    672 => X"00", 673 => X"00", 674 => X"92", 675 => X"92", 
    676 => X"54", 677 => X"54", 678 => X"38", 679 => X"FE", 
    680 => X"38", 681 => X"54", 682 => X"54", 683 => X"92", 
    684 => X"92", 685 => X"00", 686 => X"00", 687 => X"00", 
    688 => X"00", 689 => X"00", 690 => X"00", 691 => X"10", 
    692 => X"10", 693 => X"10", 694 => X"10", 695 => X"FE", 
    696 => X"10", 697 => X"10", 698 => X"10", 699 => X"10", 
    700 => X"00", 701 => X"00", 702 => X"00", 703 => X"00", 
    704 => X"00", 705 => X"00", 706 => X"00", 707 => X"00", 
    708 => X"00", 709 => X"00", 710 => X"00", 711 => X"00", 
    712 => X"00", 713 => X"08", 714 => X"08", 715 => X"10", 
    716 => X"20", 717 => X"00", 718 => X"00", 719 => X"00", 
    720 => X"00", 721 => X"00", 722 => X"00", 723 => X"00", 
    724 => X"00", 725 => X"00", 726 => X"00", 727 => X"FE", 
    728 => X"00", 729 => X"00", 730 => X"00", 731 => X"00", 
    732 => X"00", 733 => X"00", 734 => X"00", 735 => X"00", 
    736 => X"00", 737 => X"00", 738 => X"00", 739 => X"00", 
    740 => X"00", 741 => X"00", 742 => X"00", 743 => X"00", 
    744 => X"00", 745 => X"18", 746 => X"18", 747 => X"00", 
    748 => X"00", 749 => X"00", 750 => X"00", 751 => X"00", 
    752 => X"00", 753 => X"00", 754 => X"00", 755 => X"00", 
    756 => X"02", 757 => X"04", 758 => X"08", 759 => X"10", 
    760 => X"20", 761 => X"40", 762 => X"80", 763 => X"00", 
    764 => X"00", 765 => X"00", 766 => X"00", 767 => X"00", 
    768 => X"00", 769 => X"00", 770 => X"38", 771 => X"44", 
    772 => X"82", 773 => X"82", 774 => X"8A", 775 => X"92", 
    776 => X"A2", 777 => X"82", 778 => X"82", 779 => X"44", 
    780 => X"38", 781 => X"00", 782 => X"00", 783 => X"00", 
    784 => X"00", 785 => X"00", 786 => X"10", 787 => X"30", 
    788 => X"50", 789 => X"10", 790 => X"10", 791 => X"10", 
    792 => X"10", 793 => X"10", 794 => X"10", 795 => X"10", 
    796 => X"38", 797 => X"00", 798 => X"00", 799 => X"00", 
    800 => X"00", 801 => X"00", 802 => X"7C", 803 => X"82", 
    804 => X"02", 805 => X"02", 806 => X"02", 807 => X"7C", 
    808 => X"80", 809 => X"80", 810 => X"80", 811 => X"80", 
    812 => X"FE", 813 => X"00", 814 => X"00", 815 => X"00", 
    816 => X"00", 817 => X"00", 818 => X"7C", 819 => X"82", 
    820 => X"02", 821 => X"02", 822 => X"02", 823 => X"7C", 
    824 => X"02", 825 => X"02", 826 => X"02", 827 => X"82", 
    828 => X"7C", 829 => X"00", 830 => X"00", 831 => X"00", 
    832 => X"00", 833 => X"00", 834 => X"08", 835 => X"18", 
    836 => X"28", 837 => X"48", 838 => X"88", 839 => X"88", 
    840 => X"FE", 841 => X"08", 842 => X"08", 843 => X"08", 
    844 => X"1C", 845 => X"00", 846 => X"00", 847 => X"00", 
    848 => X"00", 849 => X"00", 850 => X"FE", 851 => X"80", 
    852 => X"80", 853 => X"80", 854 => X"80", 855 => X"7C", 
    856 => X"02", 857 => X"02", 858 => X"02", 859 => X"82", 
    860 => X"7C", 861 => X"00", 862 => X"00", 863 => X"00", 
    864 => X"00", 865 => X"00", 866 => X"7E", 867 => X"80", 
    868 => X"80", 869 => X"80", 870 => X"80", 871 => X"7C", 
    872 => X"82", 873 => X"82", 874 => X"82", 875 => X"82", 
    876 => X"7C", 877 => X"00", 878 => X"00", 879 => X"00", 
    880 => X"00", 881 => X"00", 882 => X"FE", 883 => X"02", 
    884 => X"02", 885 => X"04", 886 => X"08", 887 => X"10", 
    888 => X"10", 889 => X"10", 890 => X"10", 891 => X"10", 
    892 => X"38", 893 => X"00", 894 => X"00", 895 => X"00", 
    896 => X"00", 897 => X"00", 898 => X"7C", 899 => X"82", 
    900 => X"82", 901 => X"82", 902 => X"82", 903 => X"7C", 
    904 => X"82", 905 => X"82", 906 => X"82", 907 => X"82", 
    908 => X"7C", 909 => X"00", 910 => X"00", 911 => X"00", 
    912 => X"00", 913 => X"00", 914 => X"7C", 915 => X"82", 
    916 => X"82", 917 => X"82", 918 => X"82", 919 => X"7C", 
    920 => X"02", 921 => X"02", 922 => X"02", 923 => X"02", 
    924 => X"FC", 925 => X"00", 926 => X"00", 927 => X"00", 
    928 => X"00", 929 => X"00", 930 => X"00", 931 => X"00", 
    932 => X"18", 933 => X"18", 934 => X"00", 935 => X"00", 
    936 => X"00", 937 => X"18", 938 => X"18", 939 => X"00", 
    940 => X"00", 941 => X"00", 942 => X"00", 943 => X"00", 
    944 => X"00", 945 => X"00", 946 => X"00", 947 => X"00", 
    948 => X"18", 949 => X"18", 950 => X"00", 951 => X"00", 
    952 => X"00", 953 => X"08", 954 => X"08", 955 => X"10", 
    956 => X"20", 957 => X"00", 958 => X"00", 959 => X"00", 
    960 => X"00", 961 => X"00", 962 => X"00", 963 => X"00", 
    964 => X"02", 965 => X"0C", 966 => X"30", 967 => X"C0", 
    968 => X"30", 969 => X"0C", 970 => X"02", 971 => X"00", 
    972 => X"00", 973 => X"00", 974 => X"00", 975 => X"00", 
    976 => X"00", 977 => X"00", 978 => X"00", 979 => X"00", 
    980 => X"FE", 981 => X"00", 982 => X"00", 983 => X"00", 
    984 => X"00", 985 => X"00", 986 => X"FE", 987 => X"00", 
    988 => X"00", 989 => X"00", 990 => X"00", 991 => X"00", 
    992 => X"00", 993 => X"00", 994 => X"00", 995 => X"00", 
    996 => X"80", 997 => X"60", 998 => X"18", 999 => X"06", 
    1000 => X"18", 1001 => X"60", 1002 => X"80", 1003 => X"00", 
    1004 => X"00", 1005 => X"00", 1006 => X"00", 1007 => X"00", 
    1008 => X"00", 1009 => X"00", 1010 => X"38", 1011 => X"44", 
    1012 => X"82", 1013 => X"82", 1014 => X"02", 1015 => X"04", 
    1016 => X"08", 1017 => X"10", 1018 => X"10", 1019 => X"00", 
    1020 => X"10", 1021 => X"00", 1022 => X"00", 1023 => X"00", 
    1024 => X"00", 1025 => X"00", 1026 => X"38", 1027 => X"44", 
    1028 => X"82", 1029 => X"82", 1030 => X"9E", 1031 => X"A2", 
    1032 => X"A2", 1033 => X"9E", 1034 => X"80", 1035 => X"42", 
    1036 => X"3C", 1037 => X"00", 1038 => X"00", 1039 => X"00", 
    1040 => X"00", 1041 => X"00", 1042 => X"10", 1043 => X"28", 
    1044 => X"28", 1045 => X"28", 1046 => X"44", 1047 => X"7C", 
    1048 => X"44", 1049 => X"44", 1050 => X"82", 1051 => X"82", 
    1052 => X"82", 1053 => X"00", 1054 => X"00", 1055 => X"00", 
    1056 => X"00", 1057 => X"00", 1058 => X"FC", 1059 => X"82", 
    1060 => X"82", 1061 => X"82", 1062 => X"84", 1063 => X"F8", 
    1064 => X"84", 1065 => X"82", 1066 => X"82", 1067 => X"82", 
    1068 => X"FC", 1069 => X"00", 1070 => X"00", 1071 => X"00", 
    1072 => X"00", 1073 => X"00", 1074 => X"7C", 1075 => X"82", 
    1076 => X"80", 1077 => X"80", 1078 => X"80", 1079 => X"80", 
    1080 => X"80", 1081 => X"80", 1082 => X"80", 1083 => X"82", 
    1084 => X"7C", 1085 => X"00", 1086 => X"00", 1087 => X"00", 
    1088 => X"00", 1089 => X"00", 1090 => X"F0", 1091 => X"88", 
    1092 => X"84", 1093 => X"84", 1094 => X"82", 1095 => X"82", 
    1096 => X"82", 1097 => X"82", 1098 => X"84", 1099 => X"84", 
    1100 => X"F8", 1101 => X"00", 1102 => X"00", 1103 => X"00", 
    1104 => X"00", 1105 => X"00", 1106 => X"FE", 1107 => X"80", 
    1108 => X"80", 1109 => X"80", 1110 => X"80", 1111 => X"FC", 
    1112 => X"80", 1113 => X"80", 1114 => X"80", 1115 => X"80", 
    1116 => X"FE", 1117 => X"00", 1118 => X"00", 1119 => X"00", 
    1120 => X"00", 1121 => X"00", 1122 => X"FE", 1123 => X"80", 
    1124 => X"80", 1125 => X"80", 1126 => X"80", 1127 => X"FC", 
    1128 => X"80", 1129 => X"80", 1130 => X"80", 1131 => X"80", 
    1132 => X"80", 1133 => X"00", 1134 => X"00", 1135 => X"00", 
    1136 => X"00", 1137 => X"00", 1138 => X"7C", 1139 => X"82", 
    1140 => X"80", 1141 => X"80", 1142 => X"80", 1143 => X"9E", 
    1144 => X"82", 1145 => X"82", 1146 => X"82", 1147 => X"82", 
    1148 => X"7C", 1149 => X"00", 1150 => X"00", 1151 => X"00", 
    1152 => X"00", 1153 => X"00", 1154 => X"82", 1155 => X"82", 
    1156 => X"82", 1157 => X"82", 1158 => X"82", 1159 => X"7C", 
    1160 => X"82", 1161 => X"82", 1162 => X"82", 1163 => X"82", 
    1164 => X"82", 1165 => X"00", 1166 => X"00", 1167 => X"00", 
    1168 => X"00", 1169 => X"00", 1170 => X"38", 1171 => X"10", 
    1172 => X"10", 1173 => X"10", 1174 => X"10", 1175 => X"10", 
    1176 => X"10", 1177 => X"10", 1178 => X"10", 1179 => X"10", 
    1180 => X"38", 1181 => X"00", 1182 => X"00", 1183 => X"00", 
    1184 => X"00", 1185 => X"00", 1186 => X"1C", 1187 => X"08", 
    1188 => X"08", 1189 => X"08", 1190 => X"08", 1191 => X"08", 
    1192 => X"08", 1193 => X"08", 1194 => X"88", 1195 => X"88", 
    1196 => X"70", 1197 => X"00", 1198 => X"00", 1199 => X"00", 
    1200 => X"00", 1201 => X"00", 1202 => X"82", 1203 => X"82", 
    1204 => X"84", 1205 => X"84", 1206 => X"88", 1207 => X"F0", 
    1208 => X"88", 1209 => X"84", 1210 => X"84", 1211 => X"82", 
    1212 => X"82", 1213 => X"00", 1214 => X"00", 1215 => X"00", 
    1216 => X"00", 1217 => X"00", 1218 => X"80", 1219 => X"80", 
    1220 => X"80", 1221 => X"80", 1222 => X"80", 1223 => X"80", 
    1224 => X"80", 1225 => X"80", 1226 => X"80", 1227 => X"80", 
    1228 => X"FE", 1229 => X"00", 1230 => X"00", 1231 => X"00", 
    1232 => X"00", 1233 => X"00", 1234 => X"82", 1235 => X"C6", 
    1236 => X"AA", 1237 => X"AA", 1238 => X"AA", 1239 => X"92", 
    1240 => X"92", 1241 => X"82", 1242 => X"82", 1243 => X"82", 
    1244 => X"82", 1245 => X"00", 1246 => X"00", 1247 => X"00", 
    1248 => X"00", 1249 => X"00", 1250 => X"82", 1251 => X"C2", 
    1252 => X"A2", 1253 => X"A2", 1254 => X"A2", 1255 => X"92", 
    1256 => X"8A", 1257 => X"8A", 1258 => X"8A", 1259 => X"86", 
    1260 => X"82", 1261 => X"00", 1262 => X"00", 1263 => X"00", 
    1264 => X"00", 1265 => X"00", 1266 => X"7C", 1267 => X"82", 
    1268 => X"82", 1269 => X"82", 1270 => X"82", 1271 => X"82", 
    1272 => X"82", 1273 => X"82", 1274 => X"82", 1275 => X"82", 
    1276 => X"7C", 1277 => X"00", 1278 => X"00", 1279 => X"00", 
    1280 => X"00", 1281 => X"00", 1282 => X"7C", 1283 => X"82", 
    1284 => X"82", 1285 => X"82", 1286 => X"82", 1287 => X"FC", 
    1288 => X"80", 1289 => X"80", 1290 => X"80", 1291 => X"80", 
    1292 => X"80", 1293 => X"00", 1294 => X"00", 1295 => X"00", 
    1296 => X"00", 1297 => X"00", 1298 => X"7C", 1299 => X"82", 
    1300 => X"82", 1301 => X"82", 1302 => X"82", 1303 => X"82", 
    1304 => X"82", 1305 => X"B2", 1306 => X"8A", 1307 => X"84", 
    1308 => X"7A", 1309 => X"00", 1310 => X"00", 1311 => X"00", 
    1312 => X"00", 1313 => X"00", 1314 => X"7C", 1315 => X"82", 
    1316 => X"82", 1317 => X"82", 1318 => X"82", 1319 => X"FC", 
    1320 => X"A0", 1321 => X"90", 1322 => X"88", 1323 => X"84", 
    1324 => X"82", 1325 => X"00", 1326 => X"00", 1327 => X"00", 
    1328 => X"00", 1329 => X"00", 1330 => X"7C", 1331 => X"82", 
    1332 => X"80", 1333 => X"80", 1334 => X"80", 1335 => X"7C", 
    1336 => X"02", 1337 => X"02", 1338 => X"02", 1339 => X"82", 
    1340 => X"7C", 1341 => X"00", 1342 => X"00", 1343 => X"00", 
    1344 => X"00", 1345 => X"00", 1346 => X"FE", 1347 => X"92", 
    1348 => X"10", 1349 => X"10", 1350 => X"10", 1351 => X"10", 
    1352 => X"10", 1353 => X"10", 1354 => X"10", 1355 => X"10", 
    1356 => X"10", 1357 => X"00", 1358 => X"00", 1359 => X"00", 
    1360 => X"00", 1361 => X"00", 1362 => X"82", 1363 => X"82", 
    1364 => X"82", 1365 => X"82", 1366 => X"82", 1367 => X"82", 
    1368 => X"82", 1369 => X"82", 1370 => X"82", 1371 => X"82", 
    1372 => X"7C", 1373 => X"00", 1374 => X"00", 1375 => X"00", 
    1376 => X"00", 1377 => X"00", 1378 => X"82", 1379 => X"82", 
    1380 => X"82", 1381 => X"44", 1382 => X"44", 1383 => X"44", 
    1384 => X"28", 1385 => X"28", 1386 => X"28", 1387 => X"10", 
    1388 => X"10", 1389 => X"00", 1390 => X"00", 1391 => X"00", 
    1392 => X"00", 1393 => X"00", 1394 => X"82", 1395 => X"82", 
    1396 => X"82", 1397 => X"82", 1398 => X"92", 1399 => X"92", 
    1400 => X"AA", 1401 => X"AA", 1402 => X"AA", 1403 => X"C6", 
    1404 => X"82", 1405 => X"00", 1406 => X"00", 1407 => X"00", 
    1408 => X"00", 1409 => X"00", 1410 => X"82", 1411 => X"82", 
    1412 => X"44", 1413 => X"44", 1414 => X"28", 1415 => X"38", 
    1416 => X"28", 1417 => X"44", 1418 => X"44", 1419 => X"82", 
    1420 => X"82", 1421 => X"00", 1422 => X"00", 1423 => X"00", 
    1424 => X"00", 1425 => X"00", 1426 => X"82", 1427 => X"82", 
    1428 => X"44", 1429 => X"44", 1430 => X"28", 1431 => X"28", 
    1432 => X"10", 1433 => X"10", 1434 => X"10", 1435 => X"10", 
    1436 => X"10", 1437 => X"00", 1438 => X"00", 1439 => X"00", 
    1440 => X"00", 1441 => X"00", 1442 => X"FE", 1443 => X"82", 
    1444 => X"04", 1445 => X"04", 1446 => X"08", 1447 => X"38", 
    1448 => X"20", 1449 => X"40", 1450 => X"40", 1451 => X"82", 
    1452 => X"FE", 1453 => X"00", 1454 => X"00", 1455 => X"00", 
    1456 => X"00", 1457 => X"00", 1458 => X"38", 1459 => X"20", 
    1460 => X"20", 1461 => X"20", 1462 => X"20", 1463 => X"20", 
    1464 => X"20", 1465 => X"20", 1466 => X"20", 1467 => X"20", 
    1468 => X"38", 1469 => X"00", 1470 => X"00", 1471 => X"00", 
    1472 => X"00", 1473 => X"00", 1474 => X"00", 1475 => X"00", 
    1476 => X"80", 1477 => X"40", 1478 => X"20", 1479 => X"10", 
    1480 => X"08", 1481 => X"04", 1482 => X"02", 1483 => X"00", 
    1484 => X"00", 1485 => X"00", 1486 => X"00", 1487 => X"00", 
    1488 => X"00", 1489 => X"00", 1490 => X"38", 1491 => X"08", 
    1492 => X"08", 1493 => X"08", 1494 => X"08", 1495 => X"08", 
    1496 => X"08", 1497 => X"08", 1498 => X"08", 1499 => X"08", 
    1500 => X"38", 1501 => X"00", 1502 => X"00", 1503 => X"00", 
    1504 => X"00", 1505 => X"00", 1506 => X"00", 1507 => X"10", 
    1508 => X"28", 1509 => X"44", 1510 => X"82", 1511 => X"00", 
    1512 => X"00", 1513 => X"00", 1514 => X"00", 1515 => X"00", 
    1516 => X"00", 1517 => X"00", 1518 => X"00", 1519 => X"00", 
    1520 => X"00", 1521 => X"00", 1522 => X"00", 1523 => X"00", 
    1524 => X"00", 1525 => X"00", 1526 => X"00", 1527 => X"00", 
    1528 => X"00", 1529 => X"00", 1530 => X"00", 1531 => X"00", 
    1532 => X"FE", 1533 => X"00", 1534 => X"00", 1535 => X"00", 
    1536 => X"00", 1537 => X"00", 1538 => X"20", 1539 => X"20", 
    1540 => X"10", 1541 => X"10", 1542 => X"08", 1543 => X"00", 
    1544 => X"00", 1545 => X"00", 1546 => X"00", 1547 => X"00", 
    1548 => X"00", 1549 => X"00", 1550 => X"00", 1551 => X"00", 
    1552 => X"00", 1553 => X"00", 1554 => X"00", 1555 => X"00", 
    1556 => X"00", 1557 => X"00", 1558 => X"3A", 1559 => X"C6", 
    1560 => X"82", 1561 => X"82", 1562 => X"82", 1563 => X"C6", 
    1564 => X"3A", 1565 => X"00", 1566 => X"00", 1567 => X"00", 
    1568 => X"00", 1569 => X"00", 1570 => X"80", 1571 => X"80", 
    1572 => X"80", 1573 => X"80", 1574 => X"B8", 1575 => X"C6", 
    1576 => X"82", 1577 => X"82", 1578 => X"82", 1579 => X"C6", 
    1580 => X"B8", 1581 => X"00", 1582 => X"00", 1583 => X"00", 
    1584 => X"00", 1585 => X"00", 1586 => X"00", 1587 => X"00", 
    1588 => X"00", 1589 => X"00", 1590 => X"3C", 1591 => X"C2", 
    1592 => X"80", 1593 => X"80", 1594 => X"80", 1595 => X"C2", 
    1596 => X"3C", 1597 => X"00", 1598 => X"00", 1599 => X"00", 
    1600 => X"00", 1601 => X"00", 1602 => X"02", 1603 => X"02", 
    1604 => X"02", 1605 => X"02", 1606 => X"3A", 1607 => X"C6", 
    1608 => X"82", 1609 => X"82", 1610 => X"82", 1611 => X"C6", 
    1612 => X"3A", 1613 => X"00", 1614 => X"00", 1615 => X"00", 
    1616 => X"00", 1617 => X"00", 1618 => X"00", 1619 => X"00", 
    1620 => X"00", 1621 => X"00", 1622 => X"38", 1623 => X"C6", 
    1624 => X"82", 1625 => X"FC", 1626 => X"80", 1627 => X"C6", 
    1628 => X"38", 1629 => X"00", 1630 => X"00", 1631 => X"00", 
    1632 => X"00", 1633 => X"00", 1634 => X"3C", 1635 => X"42", 
    1636 => X"80", 1637 => X"80", 1638 => X"F8", 1639 => X"80", 
    1640 => X"80", 1641 => X"80", 1642 => X"80", 1643 => X"80", 
    1644 => X"80", 1645 => X"00", 1646 => X"00", 1647 => X"00", 
    1648 => X"00", 1649 => X"00", 1650 => X"00", 1651 => X"00", 
    1652 => X"00", 1653 => X"00", 1654 => X"38", 1655 => X"C6", 
    1656 => X"82", 1657 => X"7E", 1658 => X"02", 1659 => X"C6", 
    1660 => X"38", 1661 => X"00", 1662 => X"00", 1663 => X"00", 
    1664 => X"00", 1665 => X"00", 1666 => X"80", 1667 => X"80", 
    1668 => X"80", 1669 => X"80", 1670 => X"B8", 1671 => X"C6", 
    1672 => X"82", 1673 => X"82", 1674 => X"82", 1675 => X"82", 
    1676 => X"82", 1677 => X"00", 1678 => X"00", 1679 => X"00", 
    1680 => X"00", 1681 => X"00", 1682 => X"00", 1683 => X"10", 
    1684 => X"00", 1685 => X"00", 1686 => X"10", 1687 => X"10", 
    1688 => X"10", 1689 => X"10", 1690 => X"10", 1691 => X"12", 
    1692 => X"0C", 1693 => X"00", 1694 => X"00", 1695 => X"00", 
    1696 => X"00", 1697 => X"00", 1698 => X"00", 1699 => X"04", 
    1700 => X"00", 1701 => X"00", 1702 => X"04", 1703 => X"04", 
    1704 => X"04", 1705 => X"04", 1706 => X"04", 1707 => X"88", 
    1708 => X"70", 1709 => X"00", 1710 => X"00", 1711 => X"00", 
    1712 => X"00", 1713 => X"00", 1714 => X"00", 1715 => X"80", 
    1716 => X"80", 1717 => X"80", 1718 => X"86", 1719 => X"B8", 
    1720 => X"C0", 1721 => X"B0", 1722 => X"88", 1723 => X"84", 
    1724 => X"82", 1725 => X"00", 1726 => X"00", 1727 => X"00", 
    1728 => X"00", 1729 => X"00", 1730 => X"20", 1731 => X"20", 
    1732 => X"20", 1733 => X"20", 1734 => X"20", 1735 => X"20", 
    1736 => X"20", 1737 => X"20", 1738 => X"20", 1739 => X"10", 
    1740 => X"0E", 1741 => X"00", 1742 => X"00", 1743 => X"00", 
    1744 => X"00", 1745 => X"00", 1746 => X"00", 1747 => X"00", 
    1748 => X"00", 1749 => X"00", 1750 => X"AC", 1751 => X"D2", 
    1752 => X"92", 1753 => X"92", 1754 => X"92", 1755 => X"92", 
    1756 => X"92", 1757 => X"00", 1758 => X"00", 1759 => X"00", 
    1760 => X"00", 1761 => X"00", 1762 => X"00", 1763 => X"00", 
    1764 => X"00", 1765 => X"00", 1766 => X"B8", 1767 => X"C6", 
    1768 => X"82", 1769 => X"82", 1770 => X"82", 1771 => X"82", 
    1772 => X"82", 1773 => X"00", 1774 => X"00", 1775 => X"00", 
    1776 => X"00", 1777 => X"00", 1778 => X"00", 1779 => X"00", 
    1780 => X"00", 1781 => X"00", 1782 => X"38", 1783 => X"C6", 
    1784 => X"82", 1785 => X"82", 1786 => X"82", 1787 => X"C6", 
    1788 => X"38", 1789 => X"00", 1790 => X"00", 1791 => X"00", 
    1792 => X"00", 1793 => X"00", 1794 => X"00", 1795 => X"00", 
    1796 => X"00", 1797 => X"00", 1798 => X"B8", 1799 => X"C6", 
    1800 => X"82", 1801 => X"FC", 1802 => X"80", 1803 => X"80", 
    1804 => X"80", 1805 => X"00", 1806 => X"00", 1807 => X"00", 
    1808 => X"00", 1809 => X"00", 1810 => X"00", 1811 => X"00", 
    1812 => X"00", 1813 => X"00", 1814 => X"3A", 1815 => X"C6", 
    1816 => X"82", 1817 => X"7E", 1818 => X"02", 1819 => X"02", 
    1820 => X"02", 1821 => X"00", 1822 => X"00", 1823 => X"00", 
    1824 => X"00", 1825 => X"00", 1826 => X"00", 1827 => X"00", 
    1828 => X"00", 1829 => X"00", 1830 => X"B8", 1831 => X"C6", 
    1832 => X"80", 1833 => X"80", 1834 => X"80", 1835 => X"80", 
    1836 => X"80", 1837 => X"00", 1838 => X"00", 1839 => X"00", 
    1840 => X"00", 1841 => X"00", 1842 => X"00", 1843 => X"00", 
    1844 => X"00", 1845 => X"00", 1846 => X"7C", 1847 => X"82", 
    1848 => X"80", 1849 => X"7E", 1850 => X"02", 1851 => X"82", 
    1852 => X"7C", 1853 => X"00", 1854 => X"00", 1855 => X"00", 
    1856 => X"00", 1857 => X"00", 1858 => X"80", 1859 => X"80", 
    1860 => X"80", 1861 => X"80", 1862 => X"F8", 1863 => X"80", 
    1864 => X"80", 1865 => X"80", 1866 => X"80", 1867 => X"42", 
    1868 => X"3C", 1869 => X"00", 1870 => X"00", 1871 => X"00", 
    1872 => X"00", 1873 => X"00", 1874 => X"00", 1875 => X"00", 
    1876 => X"00", 1877 => X"00", 1878 => X"82", 1879 => X"82", 
    1880 => X"82", 1881 => X"82", 1882 => X"82", 1883 => X"C6", 
    1884 => X"3A", 1885 => X"00", 1886 => X"00", 1887 => X"00", 
    1888 => X"00", 1889 => X"00", 1890 => X"00", 1891 => X"00", 
    1892 => X"00", 1893 => X"00", 1894 => X"82", 1895 => X"82", 
    1896 => X"82", 1897 => X"82", 1898 => X"44", 1899 => X"28", 
    1900 => X"10", 1901 => X"00", 1902 => X"00", 1903 => X"00", 
    1904 => X"00", 1905 => X"00", 1906 => X"00", 1907 => X"00", 
    1908 => X"00", 1909 => X"00", 1910 => X"82", 1911 => X"92", 
    1912 => X"92", 1913 => X"92", 1914 => X"92", 1915 => X"92", 
    1916 => X"6C", 1917 => X"00", 1918 => X"00", 1919 => X"00", 
    1920 => X"00", 1921 => X"00", 1922 => X"00", 1923 => X"00", 
    1924 => X"00", 1925 => X"00", 1926 => X"00", 1927 => X"82", 
    1928 => X"44", 1929 => X"28", 1930 => X"38", 1931 => X"44", 
    1932 => X"82", 1933 => X"00", 1934 => X"00", 1935 => X"00", 
    1936 => X"00", 1937 => X"00", 1938 => X"00", 1939 => X"00", 
    1940 => X"00", 1941 => X"00", 1942 => X"00", 1943 => X"82", 
    1944 => X"42", 1945 => X"3C", 1946 => X"08", 1947 => X"08", 
    1948 => X"30", 1949 => X"00", 1950 => X"00", 1951 => X"00", 
    1952 => X"00", 1953 => X"00", 1954 => X"00", 1955 => X"00", 
    1956 => X"00", 1957 => X"00", 1958 => X"00", 1959 => X"FE", 
    1960 => X"04", 1961 => X"08", 1962 => X"30", 1963 => X"40", 
    1964 => X"FE", 1965 => X"00", 1966 => X"00", 1967 => X"00", 
    1968 => X"00", 1969 => X"00", 1970 => X"10", 1971 => X"20", 
    1972 => X"20", 1973 => X"20", 1974 => X"40", 1975 => X"80", 
    1976 => X"40", 1977 => X"20", 1978 => X"20", 1979 => X"20", 
    1980 => X"10", 1981 => X"00", 1982 => X"00", 1983 => X"00", 
    1984 => X"00", 1985 => X"00", 1986 => X"10", 1987 => X"10", 
    1988 => X"10", 1989 => X"10", 1990 => X"10", 1991 => X"10", 
    1992 => X"10", 1993 => X"10", 1994 => X"10", 1995 => X"10", 
    1996 => X"10", 1997 => X"00", 1998 => X"00", 1999 => X"00", 
    2000 => X"00", 2001 => X"00", 2002 => X"10", 2003 => X"08", 
    2004 => X"08", 2005 => X"08", 2006 => X"04", 2007 => X"02", 
    2008 => X"04", 2009 => X"08", 2010 => X"08", 2011 => X"08", 
    2012 => X"10", 2013 => X"00", 2014 => X"00", 2015 => X"00", 
    2016 => X"00", 2017 => X"00", 2018 => X"00", 2019 => X"00", 
    2020 => X"00", 2021 => X"00", 2022 => X"60", 2023 => X"92", 
    2024 => X"0C", 2025 => X"00", 2026 => X"00", 2027 => X"00", 
    2028 => X"00", 2029 => X"00", 2030 => X"00", 2031 => X"00", 
    2032 => X"00", 2033 => X"00", 2034 => X"00", 2035 => X"00", 
    2036 => X"00", 2037 => X"00", 2038 => X"00", 2039 => X"00", 
    2040 => X"00", 2041 => X"00", 2042 => X"00", 2043 => X"00", 
    2044 => X"00", 2045 => X"00", 2046 => X"00", 2047 => X"00", 
    others => X"00"
    -- AUTOMATICALLY GENERATED... STOP
    );
begin

  s_EN <= i_EN;
  p_rom : process (i_clock)
  begin
    if rising_edge(i_clock) then
      if s_EN = '1' then
        o_DO <= c_rom(to_integer(unsigned (i_ADDR)));
		--o_DO<= x"FF";
      end if;
    end if;
  end process p_rom;

end Behavioral;
