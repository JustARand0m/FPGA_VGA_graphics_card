-- CREATOR: Michael Braun

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TOP is
	port(
		CLK_IN: in std_logic;
	    PMOD_R, PMOD_G, PMOD_B: out std_logic_vector(3 downto 0);
	    PMOD_HS, PMOD_VS: out std_logic
	);
end TOP;

architecture BEHAV of TOP is
	-- -------------------------- components -----------------------------------
	component SYNC_GEN is
		port(
			HS, VS: out std_logic;
            ADDR: out integer;
			BLANK: out std_logic;
			PIXEL_CLK: in std_logic;
			RESET: in std_logic
		);
	end component;
	
	component BLANK_CHECK is
		port(
			R_R, R_G, R_B: out std_logic_vector(3 downto 0);
			W_R, W_G, W_B: in std_logic_vector(3 downto 0);
			BLANK: in std_logic
		);
	end component;

	component MEM_CTRL is
		port(
			R_R, R_G, R_B : out std_logic_vector(3 downto 0);
			R_ADDR: in std_logic_vector(18 downto 0);
			R_CLK: in std_logic;
			W_R, W_G, W_B : in std_logic_vector(3 downto 0);
			W_ADDR: in std_logic_vector(18 downto 0);
			W_CLK: in std_logic;
			RESET: in std_logic
		);
	end component;
	
component clk_wiz_0
port
 (-- Clock in ports
  -- Clock out ports
  clk_out1          : out    std_logic;
  clk_out2          : out    std_logic;
  -- Status and control signals
  reset             : in     std_logic;
  locked            : out    std_logic;
  clk_in1           : in     std_logic
 );
 end component;
	-- -------------------------- signals --------------------------------------
	signal BLANK: std_logic;
	-- From MEM_CTRL to BLANK_CHECK
	signal MEM_BLANK_R, MEM_BLANK_G, MEM_BLANK_B: std_logic_vector(3 downto 0);
	-- From IMG_CREATE to MEM_CTRL
	signal IMG_MEM_R, IMG_MEM_G, IMG_MEM_B: std_logic_vector(3 downto 0);
	signal W_ADDR, R_ADDR: std_logic_vector(18 downto 0);
	signal PIXEL_CLK, WRITE_CLK, SYS_CLK: std_logic;
	signal CONV_ADDR: integer;
	-- -------------------------- port maps ------------------------------------
begin
    CONV_ADDR <= to_integer(unsigned(R_ADDR));
    
	INST_SYNC_GEN: SYNC_GEN port map(
		HS        => PMOD_HS,
		VS        => PMOD_VS,
        ADDR      => CONV_ADDR,
		BLANK     => BLANK,
		PIXEL_CLK => PIXEL_CLK,
		RESET     => '0'
	);
	
	INST_BLANK_CHECK: BLANK_CHECK port map(
		R_R    => PMOD_R,
		R_G    => PMOD_G,
		R_B    => PMOD_B,
		W_R    => "0000",
		W_G    => "0000",
		W_B    => "1111",
		BLANK  => BLANK
	);

	INST_MEM_CTRL: MEM_CTRL port map(
		R_R    => MEM_BLANK_R,
		R_G    => MEM_BLANK_G,
		R_B    => MEM_BLANK_B,
		R_ADDR => R_ADDR,
		R_CLK  => PIXEL_CLK,
		W_R    => IMG_MEM_R,
		W_G    => IMG_MEM_G,
		W_B    => IMG_MEM_B,
		W_ADDR => W_ADDR,
		W_CLK  => SYS_CLK,
		RESET  => '0'
	);

	INST_CLKWIZ: clk_wiz_0 port map(
		CLK_OUT1 => SYS_CLK,
		CLK_OUT2 => PIXEL_CLK,
		reset => '0',
		CLK_IN1 => CLK_IN
	);	
end BEHAV;

